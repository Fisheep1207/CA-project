module EX_MEM
(   
    RegWrite_o,
    RegWrite_i,
    MemtoReg_o,
    MemtoReg_i,
    ALUresult_o,
    ALUresult_i,
    Readdata_o,
    Readdata_i,
    INS_11_7_o,
    INS_11_7_i,
);

endmodule