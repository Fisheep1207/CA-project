module{
    input_00_i,
    input_01_i,
    input_10_i,
    input_11_i,
    select_i,
    data_o
};
endmodule;