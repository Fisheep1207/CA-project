module ID_EX
(   
    RegWrite_o,
    RegWrite_i,
    MemtoReg_o,
    MemtoReg_i,
    MemRead_o,
    MemRead_i,
    MemWrite_o,
    MemWrite_i,
    ALUOp_o,
    ALUOp_i,
    ALUSrc_o,
    ALUSrc_i,
    Readdata1_o,
    Readdata1_i,
    Readdata2_o,
    Readdata2_i,
    Imm_o,
    Imm_i,
    ALU_o,
    ALU_i,
    INS_11_7_o,
    INS_11_7_i,
);



endmodule