module{
    Rs1_i,
    Rs2_i,
    WB_Rd_i,
    WB_RegWrite_i,
    MEM_Rd_i,
    MEM_RegWrite_i,
    ForwardA_o,
    ForwardB_o,
};

endmodule