module Hazard_Detection_Unit(
    MemRead_i,
    INS_11_7_i,
    RD1addr_i,
    RD2addr_i,
    PCWrite_o,
    Stall_o,
    No_op_o
);

endmodule